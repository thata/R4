module regfile_test;
    initial begin
        $display("hello");
    end
endmodule
