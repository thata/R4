// ALU testbench
// iverilog -g 2012 -s alu_test *.sv && ./a.out
module alu_test;
    initial begin
        $display("hello");
    end
endmodule
