module regfile(
    input logic clk, we3,
    input logic [31:0] addr1, addr2, addr3, writeData3,
    output logic [31:0] readData1, readData2
);
endmodule
