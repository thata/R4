module alu(
    input logic [31:0] in1, in2,
    input logic [2:0] funct3,
    input logic [6:0] funct7,
    output logic [31:0] result,
    output logic negative, zero
);
endmodule

